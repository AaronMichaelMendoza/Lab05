`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/24/2020 01:30:24 PM
// Design Name: 
// Module Name: addsub_test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module addsub_test();

reg a0, a1, b0, b1, m;
wire s1, s2, cout;

addsub dut(
    .a0(a0),
    .a1(a1),
    .b0(b0),
    .b1(b1),
    .m(m),
    .s1(s1),
    .s2(s2),
    .cout(cout)
    );
    
initial begin
m=0;a0=0;a1=0;b0=0;b1=0;#10;
m=0;a0=0;a1=0;b0=0;b1=1;#10;
m=0;a0=0;a1=0;b0=1;b1=0;#10;
m=0;a0=0;a1=0;b0=1;b1=1;#10;
m=0;a0=0;a1=1;b0=0;b1=0;#10;
m=0;a0=0;a1=1;b0=0;b1=1;#10;
m=0;a0=0;a1=1;b0=1;b1=0;#10;
m=0;a0=0;a1=1;b0=1;b1=1;#10;
m=0;a0=1;a1=0;b0=0;b1=0;#10;
m=0;a0=1;a1=0;b0=0;b1=1;#10;
m=0;a0=1;a1=0;b0=1;b1=0;#10;
m=0;a0=1;a1=0;b0=1;b1=1;#10;
m=0;a0=1;a1=1;b0=0;b1=0;#10;
m=0;a0=1;a1=1;b0=0;b1=1;#10;
m=0;a0=1;a1=1;b0=1;b1=0;#10;
m=0;a0=1;a1=1;b0=1;b1=1;#10;
m=1;a0=0;a1=0;b0=0;b1=0;#10;
m=1;a0=0;a1=0;b0=0;b1=1;#10;
m=1;a0=0;a1=0;b0=1;b1=0;#10;
m=1;a0=0;a1=0;b0=1;b1=1;#10;
m=1;a0=0;a1=1;b0=0;b1=0;#10;
m=1;a0=0;a1=1;b0=0;b1=1;#10;
m=1;a0=0;a1=1;b0=1;b1=0;#10;
m=1;a0=0;a1=1;b0=1;b1=1;#10;
m=1;a0=1;a1=0;b0=0;b1=0;#10;
m=1;a0=1;a1=0;b0=0;b1=1;#10;
m=1;a0=1;a1=0;b0=1;b1=0;#10;
m=1;a0=1;a1=0;b0=1;b1=1;#10;
m=1;a0=1;a1=1;b0=0;b1=0;#10;
m=1;a0=1;a1=1;b0=0;b1=1;#10;
m=1;a0=1;a1=1;b0=1;b1=0;#10;
m=1;a0=1;a1=1;b0=1;b1=1;#10;
$finish;
end

endmodule
