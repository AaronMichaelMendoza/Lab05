`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Aaron Mendoza
// 
// Create Date: 09/24/2020 01:30:24 PM
// Design Name: 
// Module Name: addsub_test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module addsub_test();

reg [1:0]a;
reg [1:0]b;
reg m;
wire cout;
wire [1:0]s;

addsub dut(
    .a(a),
    .b(b),
    .m(m),
    .s(s),
    .cout(cout)
    );
    
initial begin
m=0;a[0]=0;a[1]=0;b[0]=0;b[1]=0;#10;
m=0;a[0]=0;a[1]=0;b[0]=0;b[1]=1;#10;
m=0;a[0]=0;a[1]=0;b[0]=1;b[1]=0;#10;
m=0;a[0]=0;a[1]=0;b[0]=1;b[1]=1;#10;
m=0;a[0]=0;a[1]=1;b[0]=0;b[1]=0;#10;
m=0;a[0]=0;a[1]=1;b[0]=0;b[1]=1;#10;
m=0;a[0]=0;a[1]=1;b[0]=1;b[1]=0;#10;
m=0;a[0]=0;a[1]=1;b[0]=1;b[1]=1;#10;
m=0;a[0]=1;a[1]=0;b[0]=0;b[1]=0;#10;
m=0;a[0]=1;a[1]=0;b[0]=0;b[1]=1;#10;
m=0;a[0]=1;a[1]=0;b[0]=1;b[1]=0;#10;
m=0;a[0]=1;a[1]=0;b[0]=1;b[1]=1;#10;
m=0;a[0]=1;a[1]=1;b[0]=0;b[1]=0;#10;
m=0;a[0]=1;a[1]=1;b[0]=0;b[1]=1;#10;
m=0;a[0]=1;a[1]=1;b[0]=1;b[1]=0;#10;
m=0;a[0]=1;a[1]=1;b[0]=1;b[1]=1;#10;
m=1;a[0]=0;a[1]=0;b[0]=0;b[1]=0;#10;
m=1;a[0]=0;a[1]=0;b[0]=0;b[1]=1;#10;
m=1;a[0]=0;a[1]=0;b[0]=1;b[1]=0;#10;
m=1;a[0]=0;a[1]=0;b[0]=1;b[1]=1;#10;
m=1;a[0]=0;a[1]=1;b[0]=0;b[1]=0;#10;
m=1;a[0]=0;a[1]=1;b[0]=0;b[1]=1;#10;
m=1;a[0]=0;a[1]=1;b[0]=1;b[1]=0;#10;
m=1;a[0]=0;a[1]=1;b[0]=1;b[1]=1;#10;
m=1;a[0]=1;a[1]=0;b[0]=0;b[1]=0;#10;
m=1;a[0]=1;a[1]=0;b[0]=0;b[1]=1;#10;
m=1;a[0]=1;a[1]=0;b[0]=1;b[1]=0;#10;
m=1;a[0]=1;a[1]=0;b[0]=1;b[1]=1;#10;
m=1;a[0]=1;a[1]=1;b[0]=0;b[1]=0;#10;
m=1;a[0]=1;a[1]=1;b[0]=0;b[1]=1;#10;
m=1;a[0]=1;a[1]=1;b[0]=1;b[1]=0;#10;
m=1;a[0]=1;a[1]=1;b[0]=1;b[1]=1;#10;
$finish;
end

endmodule
